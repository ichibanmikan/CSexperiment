library ieee;
use ieee.std_logic_1164.all;  --�����ͳ����

entity rom is
    port(   a4, a3, a2, a1, a0: in std_logic; --5���������΢��ַ����
            d: out std_logic_vector(28 downto 1)); --28λ������������������28λ΢ָ�����
end rom; --����ʵ��˿�

architecture rom of rom is
    signal temp: std_logic_vector(28 downto 1);
    signal a:std_logic_vector(4 downto 0);
begin
    a<=a4&a3&a2&a1&a0; --�������5����΢��ַ����ϲ���5λ������
    temp<=
		"1010111100000000000000000001"   when a="00000"else
		"1111111000001000000000000010"   when a="00001"else
		"1001111100000100000001101000"   when a="00010"else
		"1111111000001000000000010101"   when a="01001"else
		"1001111100001000000001010110"   when a="10101"else
		"1001111110000000000001000001"   when a="10110"else
		"1111111000001000000000010111"   when a="01010"else
		"1001111100001000000001011000"   when a="10111"else
		"1001101100000000000010000001"   when a="11000"else
		"1111111000001000000000011001"   when a="01011"else
		"1001111100001000000001011010"   when a="11001"else
		"1001111100000000000001000001"   when a="11010"else
		"1001101100010000000000011011"   when a="01100"else
		"1001110110000010000000000001"   when a="11011"else
		"1111111000001000000000011100"   when a="01101"else
		"1011111100000000000001000001"   when a="11100"else
		"1111111000001000000000000011"   when a="01110"else
		"1001111100001000000001000100"   when a="00011"else
		"1001111100100000000001000101"   when a="00100"else
		"1001101100010000000000000110"   when a="00101"else
		"1001110110000001100100000001"   when a="00110"else
		"1111111000001000000000011101"   when a="01111"else
		"1001111100001000000001011110"   when a="11101"else
		"1001111100100000000001011111"   when a="11110"else
		"1001101100010000000000000111"   when a="11111"else
		"1001110110000000101100000001"   when a="00111"else
		"1010111100000000000000010001"   when a="10000"else
		"1111111000001000000000010010"   when a="10001"else
		"1000111100000000000010010001"   when a="10010"else
		"1010111100000000000000010011"   when a="01000"else
		"1111111000001000000000010100"   when a="10011"else
		"1001111100000000000001010011"   when a="10100"; --�������
    d <= temp;
end rom;